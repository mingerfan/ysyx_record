module top();
endmodule

